
`define frac 12
`define exp 8
