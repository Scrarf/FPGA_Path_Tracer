module 16bit_LZC (
	input clk,

);

endmodule