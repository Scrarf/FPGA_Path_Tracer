`include "src/arithmetic_cores/definitions.vh"

/*
Inputs are unpacked arrays.
Only works for Normalized non-special case numbers.
Needs propper zero handling at least.

The module is pipelined.
*/

module add (
	input wire clk,
	input u_float a,
	input u_float b,
	output u_float c
);

reg [`exp:0] exp_diff, exp_diff_abs, exp_greater, exp_greater_dl, exp_greater_dl2, exp_greater_dl3, exp_greater_dl4, exp_greater_dl5, exp_greater_dl6;
reg [`exp:0] exp_greater_normalized, exp_greater_normalized_dl, exp_greater_normalized_dl2;
reg sign_xor, sign_xor_dl, sign_xor_dl2;
reg sign_c, sign_c_dl, sign_c_dl2, sign_c_dl3, sign_c_dl4, sign_c_dl5, sign_c_dl6, sign_c_dl7, sign_c_dl8, sign_c_dl9;
reg [`frac:0] frac_to_be_shifted, frac_to_be_shifted_dl, frac_to_be_bypassed, frac_to_be_bypassed_dl, frac_to_be_bypassed_dl2, frac_to_be_bypassed_dl3;
reg [(`frac*2)+1:0] frac_shifted;
reg [(`frac*2)+3:0] frac_shifted_inverted;
reg [(`frac*2)+3:0] frac_combined, frac_combined_abs, frac_combined_abs_dl;
reg [`frac:0] frac_normalized_trunk, frac_normalized;
reg [`frac+1:0] frac_normalized_trunk_rounded;

reg round_up, round, guard, sticky;

sixteen_bit_lzc LZC(.clk(clk), .array(frac_combined_abs[(`frac*2)+3:(`frac*2)-12]), .value(lzc));
reg [3:0] lzc;

wire exp_comparison = $signed(a.exp) > $signed(b.exp);
//11 pipeline stages
always @(posedge clk) begin
	/*===========================================================*/
	exp_diff <= a.exp - b.exp;
	exp_greater <= exp_comparison ? a.exp : b.exp;
	
	frac_to_be_shifted <= exp_comparison ? b.frac : a.frac;
	frac_to_be_bypassed <= exp_comparison ? a.frac : b.frac;

	sign_xor <= a.sign ^ b.sign;
	sign_c <= (a.exp == b.exp) ? ((a.frac > b.frac) ? a.sign : b.sign) : (exp_comparison ? a.sign : b.sign);

	/*===========================================================*/
	sign_xor_dl <= sign_xor;
	sign_c_dl <= sign_c;

	exp_greater_dl <= exp_greater;
	exp_diff_abs <= exp_diff[`exp] ? (~exp_diff + 1'b1) : exp_diff;

	frac_to_be_shifted_dl <= frac_to_be_shifted;
	frac_to_be_bypassed_dl <= frac_to_be_bypassed;

	/*===========================================================*/
	sign_xor_dl2 <= sign_xor_dl;

	exp_greater_dl2 <= exp_greater_dl;

	frac_shifted <= {frac_to_be_shifted_dl, `frac'b0, 1'b0} >> exp_diff_abs; //2x size of frac_to_be_shifted
	frac_to_be_bypassed_dl2 <= frac_to_be_bypassed_dl;

	sign_c_dl2 <= sign_c_dl;

	/*===========================================================*/
	exp_greater_dl3 <= exp_greater_dl2;

	frac_shifted_inverted <= sign_xor_dl2 ? (~({2'b0, frac_shifted}) + 1'b1) : {2'b0, frac_shifted};
	frac_to_be_bypassed_dl3 <= frac_to_be_bypassed_dl2;

	sign_c_dl3 <= sign_c_dl2;

	/*===========================================================*/
	exp_greater_dl4 <= exp_greater_dl3;

	frac_combined <= {2'b0, frac_to_be_bypassed_dl3, `frac'b0, 1'b0} + frac_shifted_inverted;

	sign_c_dl4 <= sign_c_dl3;

	/*===========================================================*/
	exp_greater_dl5 <= exp_greater_dl4;

	frac_combined_abs <= frac_combined[(`frac*2)+3] ? (~frac_combined + 1'b1) : frac_combined;

	sign_c_dl5 <= sign_c_dl4;

	/*===========================================================*/
	exp_greater_dl6 <= exp_greater_dl5;
	//LZC here
	frac_combined_abs_dl <= frac_combined_abs;

	sign_c_dl6 <= sign_c_dl5;

	/*===========================================================*/
	exp_greater_normalized <= (exp_greater_dl6 - {5'b0, lzc}) + 2;
	
	frac_normalized <= {frac_combined_abs_dl << lzc}[(`frac*2)+3:(`frac+3)]; //UNUSED SIGNAL WARNING

	guard <= {(frac_combined_abs_dl << lzc)}[`frac+2];
	round <= {(frac_combined_abs_dl << lzc)}[`frac+1];
	sticky <= |{(frac_combined_abs_dl << lzc)}[`frac:0];

	sign_c_dl7 <= sign_c_dl6;

	/*===========================================================*/
	exp_greater_normalized_dl <= exp_greater_normalized;

	frac_normalized_trunk <= frac_normalized;

	sign_c_dl8 <= sign_c_dl7;

	round_up <= guard & (round | sticky | frac_normalized[0]);
	/*===========================================================*/
	exp_greater_normalized_dl2 <= exp_greater_normalized_dl;

	frac_normalized_trunk_rounded <= {1'b0, frac_normalized_trunk} + {{(`frac){1'b0}}, round_up};

	sign_c_dl9 <= sign_c_dl8;

	/*===========================================================*/
	c.sign <= sign_c_dl9;
	//c.sign <= 1;

	//{1'b0, c.frac} <= frac_normalized_trunk_rounded >> frac_normalized_trunk_rounded[`frac+1];
	c.frac <= {frac_normalized_trunk_rounded >> frac_normalized_trunk_rounded[`frac+1]}[12:0];

	c.exp <= exp_greater_normalized_dl2 + {`exp'b0, frac_normalized_trunk_rounded[`frac+1]};


end

endmodule

/*
NEXTPNR REPORT:

Max frequency: 199.64 MHz.

Info: Device utilisation:
Info:             TRELLIS_IO:      70/    365    19%
Info:                   DCCA:       1/     56     1%
Info:                 DP16KD:       0/    208     0%
Info:             MULT18X18D:       0/    156     0%
Info:                 ALU54B:       0/     78     0%
Info:                EHXPLLL:       0/      4     0%
Info:                EXTREFB:       0/      2     0%
Info:                   DCUA:       0/      2     0%
Info:              PCSCLKDIV:       0/      2     0%
Info:                IOLOGIC:       0/    224     0%
Info:               SIOLOGIC:       0/    141     0%
Info:                    GSR:       0/      1     0%
Info:                  JTAGG:       0/      1     0%
Info:                   OSCG:       0/      1     0%
Info:                  SEDGA:       0/      1     0%
Info:                    DTR:       0/      1     0%
Info:                USRMCLK:       0/      1     0%
Info:                CLKDIVF:       0/      4     0%
Info:              ECLKSYNCB:       0/     10     0%
Info:                DLLDELD:       0/      8     0%
Info:                 DDRDLL:       0/      4     0%
Info:                DQSBUFM:       0/     14     0%
Info:        TRELLIS_ECLKBUF:       0/      8     0%
Info:           ECLKBRIDGECS:       0/      2     0%
Info:                   DCSC:       0/      2     0%
Info:             TRELLIS_FF:     399/  83640     0%
Info:           TRELLIS_COMB:     765/  83640     0%
Info:           TRELLIS_RAMW:       0/  10455     0%

*/
